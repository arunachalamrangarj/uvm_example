`define HDR "**********************************************"
`define HDR_LINE  "This is my Hello World test"
`define PREFIX "My simple test"